`timescale 1ps / 1ps

module Address_decoder ();



endmodule
