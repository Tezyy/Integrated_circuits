*Mem_cell
*Logic gates (V1 untested 19_10)


.include gpdk90nm_tt.cir


*Logic gates (V1 untested 19_10)


*________________________________________________

*NOT gate 

.subckt 1inNOT in1 out1 Vdd gnd
xMp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xMn1 out1 in1 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________

*NAND gates

.subckt 2inNAND in1 in2 out1 Vdd gnd
xmp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp2 Vdd in2 out1 Vdd pmos1v L=Lpmos W=Wpmos

xmn1 out1 in1 2 gnd nmos1v L=L1 W=W1
xmn2 2 in2 gnd gnd nmos1v L=L1 W=W1
.ends

.subckt 3inNAND in1 in2 in3 out1 Vdd gnd
xmp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp2 Vdd in2 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp3 Vdd in3 out1 Vdd pmos1v L=Lpmos W=Wpmos

xmn1 out1 in1 2 gnd nmos1v L=L1 W=W1
xmn2 2 in2 3 gnd nmos1v L=L1 W=W1
xmn3 3 in3 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________

*AND gates

.subckt 2inAND in1 in2 out1 Vdd gnd
xNAND1 in1 in2 temp Vdd gnd 2inNAND
xNOT1 temp out1 Vdd gnd 1inNOT
.ends

.subckt 3inAND in1 in2 in3 out1 Vdd gnd
xNAND1 in1 in2 in3 temp Vdd gnd 3inNAND
xNOT1 temp out1 Vdd gnd 1inNOT
.ends

*________________________________________________

*NOR gate

.subckt 2inNOR in1 in2 out1 Vdd gnd
xmp1 Vdd in1 dp2 Vdd pmos1v L=L1 W=W1
xmp2 dp2 in2 out1 Vdd pmos1v L=L1 W=W1

xmn1 out1 in1 gnd gnd nmos1v L=L1 W=W1
xmn2 out1 in2 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________


*paramètres
*Transistor dimensions: 100nm < W < 1500nm and 100nm < L < 300nm
* 0.4 < Vdd < 1
.param Vdd=1
.param L1=100n
.param W1=300n
.param Lpmos=100n
.param Wpmos=750n




.subckt SR_latch in1 in2 out1 Vdd gnd
xNAND1 in1 not_out out1 Vdd gnd 2inNAND
xNAND2 out1 in2 not_out Vdd gnd 2inNAND
.ends

.subckt Bitcell select input rw out_bitcell out_SRlatch Vdd gnd

xNAND1 select input rw outNAND1 Vdd gnd 3inNAND
xNAND2 select outNAND1 rw outNAND2 Vdd gnd 3inNAND

xNOT2 rw not_rw Vdd gnd 1inNOT

xAND3 not_rw out_SRLATCH select out_bitcell Vdd gnd 3inAND

xSRLATCH outNAND1 outNAND2 out_SRLATCH Vdd gnd SR_latch

.ends


*______________________________________________

*FOR THE TESTS : COPY & PASTE THE SPICE CODE FROM
*THE WANTED FILES

V1 1 0 dc Vdd
Vinp in 0 PULSE(0 Vdd 0ns 0.1ns 0.1ns 10ns 100ns)
Vsel sel 0 PULSE(0 Vdd 0ns 0.1ns 0.1ns 100ns 100ns)
Vrw rw 0 PULSE(0 Vdd 25ns 0.1ns 0.1ns 10ns 20ns)


*Testing read/write time
xBitcell sel in rw YYYY_cell YYYY_latch 1 0 bitcell
.plot v(in) v(sel) v(rw) v(YYYY_cell) v(YYYY_latch)
.plot v(YYYY_cell) v(YYYY_latch)

.plot i(V1)


*_______________________________________________________



*_______________________________________________________