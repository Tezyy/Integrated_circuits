*Mem_cell
*Logic gates (V1 untested 19_10)


.include gpdk90nm_tt.cir


*Logic gates (V1 untested 19_10)


*________________________________________________

*NOT gate 

.subckt 1inNOT in1 out1 Vdd gnd
xMp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xMn1 out1 in1 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________

*NAND gates

.subckt 2inNAND in1 in2 out1 Vdd gnd
xmp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp2 Vdd in2 out1 Vdd pmos1v L=Lpmos W=Wpmos

xmn1 out1 in1 2 gnd nmos1v L=L1 W=W1
xmn2 2 in2 gnd gnd nmos1v L=L1 W=W1
.ends

.subckt 3inNAND in1 in2 in3 out1 Vdd gnd
xmp1 Vdd in1 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp2 Vdd in2 out1 Vdd pmos1v L=Lpmos W=Wpmos
xmp3 Vdd in3 out1 Vdd pmos1v L=Lpmos W=Wpmos

xmn1 out1 in1 2 gnd nmos1v L=L1 W=W1
xmn2 2 in2 3 gnd nmos1v L=L1 W=W1
xmn3 3 in3 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________

*AND gates

.subckt 2inAND in1 in2 out1 Vdd gnd
xNAND1 in1 in2 temp Vdd gnd 2inNAND
xNOT1 temp out1 Vdd gnd 1inNOT
.ends

.subckt 3inAND in1 in2 in3 out1 Vdd gnd
xNAND1 in1 in2 in3 temp Vdd gnd 3inNAND
xNOT1 temp out1 Vdd gnd 1inNOT
.ends

*________________________________________________

*NOR gate

.subckt 2inNOR in1 in2 out1 Vdd gnd
xmp1 Vdd in1 dp2 Vdd pmos1v L=L1 W=W1
xmp2 dp2 in2 out1 Vdd pmos1v L=L1 W=W1

xmn1 out1 in1 gnd gnd nmos1v L=L1 W=W1
xmn2 out1 in2 gnd gnd nmos1v L=L1 W=W1
.ends

*________________________________________________


*paramètres
*  Transistor dimensions: 100nm < W < 1500nm and 100nm < L < 300nm
.param Vdd=1
.param L1=200n
.param W1=600n
.param Lpmos=200n
.param Wpmos=1500n




.subckt SR_latch in1 in2 out1 Vdd gnd
xNAND1 in1 not_out out1 Vdd gnd 2inNAND
xNAND2 out1 in2 not_out Vdd gnd 2inNAND
.ends

.subckt bitcell select input rw out_bitcell out_SRlatch Vdd gnd

xNAND1 select input rw outNAND1 Vdd gnd 3inNAND
xNAND2 select outNAND1 rw outNAND2 Vdd gnd 3inNAND

xNOT2 rw not_rw Vdd gnd 1inNOT

xAND3 not_rw out_SRLATCH select out_bitcell Vdd gnd 3inAND

xSRLATCH outNAND1 outNAND2 out_SRLATCH Vdd gnd SR_latch

.ends


*______________________________________________

*Test signals
V1 1 0 dc Vdd
Vinp in 0 PULSE(0 Vdd 35ns 0.1ns 0.1ns 10ns 50ns)
Vsel sel 0 PULSE(0 Vdd 15ns 0.1ns 0.1ns 5ns 10ns)
Vrw rw 0 PULSE(0 Vdd 10ns 0.1ns 0.1ns 10ns 20ns)

*Vinp in 0 PULSE(0 Vdd 35ns 0.1ns 0.1ns 25ns 50ns)
*Vsel sel 0 PULSE(0 Vdd 15ns 0.1ns 0.1ns 25ns 50ns)
*Vrw rw 0 PULSE(0 Vdd 10ns 0.1ns 0.1ns 20ns 40ns)

*Testing read/write time
xBitcell sel in rw YYYY_cell YYYY_latch 1 0 bitcell
.plot v(in) v(sel) v(rw) v(YYYY_cell) v(YYYY_latch)
*.plot i(v1)

*leakage measurement
*xBitcell 0 1 1 YYYY_cell YYYY_latch 1 0 SRbitcell
*.op xBitcell


*_______________________________________________________


*TEST LOGICAL GATES 
*NOT : ok NAND_3IN 
Vdd voltage 0 dc Vdd
Vin1 in1 0 PULSE(0 Vdd 0 1n 1n 10n 20n)
Vin2 in2 0 PULSE(0 Vdd 0 1n 1n 20n 40n)
Vin3 in3 0 PULSE(0 Vdd 0 1n 1n 40n 80n)


* Test 1-input NOT gate
xNOT_test in1 out_not voltage 0 1inNOT
* Test 2-input AND gate
xAND2_test in1 in2 out_and2 voltage 0 2inAND
* Test 3-input AND gate
xAND3_test in1 in2 in3 out_and3 voltage 0 3inAND
* Test 2-input NOR gate
xNOR2_test in1 in2 out_nor2 voltage 0 2inNOR
* Test 3-input NAND gate
xNAND3_test in1 in2 in3 out_nand3 voltage 0 3inNAND

* Test 2-input NAND gate
xNAND2_test in1 in2 out_nand2 voltage 0 2inNAND

* Test SRLATCH gate
xlatch in1 in2 out_latch voltage 0 SR_latch

xNAND1 in1 in2 in3 outNAND1 voltage 0 3inNAND
xNAND2 outNAND1 in1 in2 outNAND2 voltage 0 3inNAND

